--------------------------------------------------------------------------------
-- Company: 		Binghamton University
-- Engineer:		Carl Betcher
--
-- Create Date:   21:31:25 04/16/2011
-- Design Name:   Lab 7C Testbench
-- Module Name:   Test_Lab7C.vhd
-- Project Name:  Lab7
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Lab7C_top_level
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
--	   04/04/2015 - Modified the process to verify the nrz_out data matches
--						 the Machester data generated by the stimulus process
--					  - Generalized to work for different system clock speeds
-- Additional Comments:
--
-- Notes: 
-- Run this simulation for 40 us (Papilio) or 25 us (Basys2)
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY Test_Lab7C IS
END Test_Lab7C;
 
ARCHITECTURE behavior OF Test_Lab7C IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Lab7C_top_level
	 GENERIC (debounceDELAY : integer := 640000); 
    PORT(
         manin : IN  std_logic;
         manout : OUT  std_logic;
         dclk_in : IN  std_logic;
         frame_in : IN  std_logic;
         nrz_in : IN  std_logic;
			dclk_out : OUT STD_LOGIC;
			frame_out : OUT STD_LOGIC;
         nrz_out : OUT  std_logic;
         mclk : IN  std_logic;
         rst : IN  std_logic
        );
    END COMPONENT;
    
   --Inputs
   signal manin : std_logic := '0';
   signal dclk_in : std_logic := '0';
   signal frame_in : std_logic := '0';
   signal nrz_in : std_logic := '0';
   signal mclk : std_logic := '0';
   signal rst : std_logic := '0';

 	--Outputs
   signal manout : std_logic;
   signal dclk_out : std_logic;
   signal frame_out : std_logic;
   signal nrz_out : std_logic;

   -- Clock period definitions
--	constant mclk_period : time := 20 ns;    -- Basys2
	constant mclk_period : time := 31.25 ns; -- Papilio

	constant txdata_period : time := 32*mclk_period;
									-- period of each data bit sent
									-- is the period of 32 system clocks

	-- Test Data
	type test_array_type is array (natural range <>) of std_logic_vector(7 downto 0);	
	constant test_data : test_array_type :=
		(
			("10101010"),   -- Preamble
			("10101011"),   -- Start Frame Delimiter (SFD)
			("00001111"),   -- Data
			("00110011")    -- Data
		);
	
	signal data_byte : std_logic_vector(7 downto 0) := (others => '0');	

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Lab7C_top_level 
	GENERIC MAP ( debounceDELAY => 3 )  
	PORT MAP (
          manin => manin,
          manout => manout,
          dclk_in => dclk_in,
          frame_in => frame_in,
          nrz_in => nrz_in,
			 dclk_out => dclk_out,
			 frame_out => frame_out,
          nrz_out => nrz_out,
          mclk => mclk,
          rst => rst
        );

   -- Clock process definitions
   mclk_process :process
   begin
		mclk <= '0';
		wait for mclk_period/2;
		mclk <= '1';
		wait for mclk_period/2;
   end process;
 
 	-- External connections
	manin <= manout;

   -- Results Checking Process
	-- This process is separate from the stimulus process,
	-- waits for the rising edge of frame_out and checks
	-- that the NRZ_out data matches the Manchester data 
	-- that was sent by the stimulus process
   check_proc: process
		variable error_flag : std_logic := '0';
	begin
		wait until rising_edge(frame_out);
		error_flag := '0';
		report "testing for bad NRZ bit values" severity NOTE;
		for j in 0 to 3 loop
			data_byte <=test_data(j);
			for k in 7 downto 0 loop
				wait until rising_edge(dclk_out);
				-- test that decoded NRZ equals encoded data bit
				if nrz_out /= data_byte(k) then error_flag := '1'; end if;
				assert nrz_out = data_byte(k)
					report "NRZ_OUT does not equal Manchester data bit" 
					severity ERROR;
				wait until falling_edge(dclk_out);
			end loop;
		end loop;
		if error_flag = '0' then report "NO ERRORS FOUND" severity NOTE; end if;
   end process;
	
	-- Stimulus process
   stim_proc: process
	
	procedure tx_data_byte (data: in std_logic_vector(7 downto 0)) is
	begin
		for I in 7 downto 0 loop
			nrz_in <= data(I);
			wait for txdata_period/2;
			dclk_in <= '1';
			wait for txdata_period/2;
			dclk_in <= '0';
		end loop;
	end procedure;
	
   begin	
		-- initialization
		nrz_in <= '0';
		dclk_in <= '0';
		frame_in <= '0';
      -- generate reset
		rst <= '0';
      wait for mclk_period*5;	
		rst <= '1';
      wait for mclk_period*5;	
		rst <= '0';

      wait for 1.8 us;

      -- insert stimulus here 
		-- generate nrz data to be transmitted
		frame_in <= '1';
		for i in test_data'range loop
			tx_data_byte(test_data(i));   -- transmit a data byte
		end loop;
		frame_in <= '0';
		nrz_in <= '0';

      wait;
   end process;
	
END;
