--------------------------------------------------------------------------------
-- Company: 		Binghamton University
-- Engineer:		Carl Betcher
--
-- Create Date:   17:48:34 04/17/2011
-- Design Name:   Lab 7C Testbench for Manchester Decoder Only
-- Module Name:   Test_Lab7C_md.vhd
-- Project Name:  Lab7
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: manchdecoder
-- 
-- Dependencies:
-- 
-- Revisions:
-- Revision 0.01 - File Created
--	   04/04/2015 - Added separate process to verify the nrz_out data matches
--						 the Machester data generated by the stimulus process
--					  - Modified the stimulus procedure to generate the entire
--						 frame instead of a byte of data
--					  - Generalized to work for different system clock speeds
-- Additional Comments:
--
-- Notes: 
-- Run this simulation for 120 usec (Papilio) or 80 usec (Basys2)
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY Test_Lab7C_md IS
END Test_Lab7C_md;
 
ARCHITECTURE behavior OF Test_Lab7C_md IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT manchdecoder
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         manin : IN  std_logic;
         dclk_out : OUT  std_logic;
         frame_out : OUT  std_logic;
         nrz_out : OUT  std_logic
        );
    END COMPONENT;
    
   --Inputs
   signal rst : std_logic := '0';
   signal clk : std_logic := '0';
   signal manin : std_logic := '0';

 	--Outputs
   signal dclk_out : std_logic;
   signal frame_out : std_logic;
   signal nrz_out : std_logic;

   -- Clock period definitions
--	constant clk_period : time := 20 ns;    -- Basys2
	constant clk_period : time := 31.25 ns; -- Papilio

	shared variable man_clk_period : time := 32*clk_period;
									-- period of each data bit sent
									-- is the period of 32 system clocks
									-- shared variable allows testing of the
									-- affects of clock frequency variations

	-- Clock to establish Manchester signal timing
	signal tb_man_clk : std_logic;
	
	-- Test data - four bytes of data used in each frame
	type test_array_type is array (natural range <>) of std_logic_vector(7 downto 0);
	constant TEST_ARRAY: test_array_type :=
		(
			("10101010"),
			("10101011"),
			("00001111"),
			("00110011")
		);

	signal check_NRZ : std_logic := '0';

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: manchdecoder PORT MAP (
          rst => rst,
          clk => clk,
          manin => manin,
          dclk_out => dclk_out,
          frame_out => frame_out,
          nrz_out => nrz_out
        );

   -- Clock process definitions
	-- System Clock
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   -- Manchester Clock
	man_clk_process :process
   begin
		tb_man_clk <= '0';
		wait for man_clk_period/2;
		tb_man_clk <= '1';
		wait for man_clk_period/2;
   end process;
 
   -- Results Checking Process
	-- This process is separate from the stimulus process,
	-- waits for the rising edge of frame_out and checks
	-- that the NRZ_out data matches the Manchester data 
	-- that was sent by the stimulus process
   check_proc: process
		variable byte : std_logic_vector(7 downto 0);
		variable error_flag : std_logic := '0';
	begin
		for i in 0 to 2 loop
			wait until rising_edge(frame_out);
			error_flag := '0';
			report "testing for bad NRZ bit values" severity NOTE;
			for j in 0 to 3 loop
				byte := TEST_ARRAY(j);
				for k in 7 downto 0 loop
					wait until rising_edge(dclk_out);
					-- test that decoded NRZ equals encoded data bit
					check_NRZ <= '1';
					if nrz_out /= byte(k) then error_flag := '1'; end if;
					assert nrz_out = byte(k)
						report "NRZ_OUT does not equal Manchester data bit" 
						severity ERROR;
					wait until falling_edge(dclk_out);
					check_NRZ <= '0';
				end loop;
			end loop;
			if error_flag = '0' then report "NO ERRORS FOUND" severity NOTE; end if;
		end loop;
   end process;
	
   -- Stimulus Process
   stim_proc: process
	
	-- procedure to generate a frame of Manchester data on manin
	-- using data from TEST_ARRAY
	procedure manch_frame(TEST_ARRAY : in test_array_type) is
		variable data : std_logic_vector(7 downto 0);
	begin
		for i in TEST_ARRAY'range loop
			data := TEST_ARRAY(i);
			for j in data'range loop
				-- encode data bit
				wait until falling_edge(tb_man_clk);
				if data(j) = '1' then manin <= '0'; else manin <= '1'; end if;	
				wait until rising_edge(tb_man_clk);
				if data(j) = '1' then manin <= '1'; else manin <= '0'; end if;	
			end loop;	
		end loop;		
	end procedure;
	
   begin
		manin <= '0';
		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		rst <= '0';
      wait for 100 ns;	
		rst <= '1';
      wait for 100 ns;	
		rst <= '0';

      wait for 4.7 us;
		
      -- insert stimulus here
		-- generate Manchester data on manin using nominal clock period
		report "Manchester clock period = nominal value" severity NOTE;
		manch_frame(TEST_ARRAY);
		wait until falling_edge (tb_man_clk);
		manin <= '0';
		wait for 2.5 us;

		-- generate Manchester data on manin using nominal clock period - 10%
		report "Manchester clock period = 10% low" severity NOTE;
		man_clk_period := 32*clk_period-(32*clk_period*0.10); -- clock period is 10% low
		wait for 2.5 us;
		manch_frame(TEST_ARRAY);
		wait until falling_edge (tb_man_clk);
		manin <= '0';
		wait for 2.5 us;

		-- generate Manchester data on manin using nominal clock period + 10%
		report "Manchester clock period = 10% high" severity NOTE;
		man_clk_period := 32*clk_period*1.10; -- clock period is 10% high
		wait for 2.5 us;
		manch_frame(TEST_ARRAY);
		wait until falling_edge (tb_man_clk);
		manin <= '0';

      wait;
   end process;

END;